
module lab7_soc (
	clk_clk,
	led_wire_export,
	sdram_clk_clk,
	sdram_wire_addr,
	sdram_wire_ba,
	sdram_wire_cas_n,
	sdram_wire_cke,
	sdram_wire_cs_n,
	sdram_wire_dq,
	sdram_wire_dqm,
	sdram_wire_ras_n,
	sdram_wire_we_n,
	sw_wire_export,
	acc_wire_export,
	reset_reset_n,
	reset_wire_export);	

	input		clk_clk;
	output	[7:0]	led_wire_export;
	output		sdram_clk_clk;
	output	[12:0]	sdram_wire_addr;
	output		sdram_wire_ba;
	output		sdram_wire_cas_n;
	output		sdram_wire_cke;
	output	[1:0]	sdram_wire_cs_n;
	inout	[31:0]	sdram_wire_dq;
	output	[3:0]	sdram_wire_dqm;
	output		sdram_wire_ras_n;
	output		sdram_wire_we_n;
	input	[7:0]	sw_wire_export;
	input		acc_wire_export;
	input		reset_reset_n;
	input		reset_wire_export;
endmodule
